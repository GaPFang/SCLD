// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 32-bit"
// VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
// CREATED		"Wed Dec 28 16:57:18 2022"

module DataReg(
	rst_n,
	clk,
	A,
	Q
);


input wire	rst_n;
input wire	clk;
input wire	[3:0] A;
output wire	[3:0] Q;

wire	[3:0] Q_ALTERA_SYNTHESIZED;





DFF_1	b2v_inst(
	.CLK(clk),
	.D(A[3]),
	
	.ClrN(rst_n),
	
	.Q(Q_ALTERA_SYNTHESIZED[3]));


DFF_1	b2v_inst1(
	.CLK(clk),
	.D(A[2]),
	
	.ClrN(rst_n),
	
	.Q(Q_ALTERA_SYNTHESIZED[2]));


DFF_1	b2v_inst2(
	.CLK(clk),
	.D(A[1]),
	
	.ClrN(rst_n),
	
	.Q(Q_ALTERA_SYNTHESIZED[1]));


DFF_1	b2v_inst5(
	.CLK(clk),
	.D(A[0]),
	
	.ClrN(rst_n),
	
	.Q(Q_ALTERA_SYNTHESIZED[0]));

assign	Q = Q_ALTERA_SYNTHESIZED;

endmodule
