library verilog;
use verilog.vl_types.all;
entity FS_vlg_vec_tst is
end FS_vlg_vec_tst;
